library verilog;
use verilog.vl_types.all;
entity newspaper_test is
end newspaper_test;
