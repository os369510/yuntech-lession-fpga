library verilog;
use verilog.vl_types.all;
entity adder_8bit_tb1 is
end adder_8bit_tb1;
