library verilog;
use verilog.vl_types.all;
entity BCD_adder_test is
end BCD_adder_test;
